library verilog;
use verilog.vl_types.all;
entity displayController_vlg_vec_tst is
end displayController_vlg_vec_tst;
