library verilog;
use verilog.vl_types.all;
entity displayController_vlg_check_tst is
    port(
        DisplayOut      : in     vl_logic_vector(7 downto 0);
        sampler_rx      : in     vl_logic
    );
end displayController_vlg_check_tst;
