library verilog;
use verilog.vl_types.all;
entity eight_bit_reg_shift_r_vlg_vec_tst is
end eight_bit_reg_shift_r_vlg_vec_tst;
